package piso_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // Import sub-packages
    import piso_sequences_pkg::*;
    import piso_agent_pkg::*;
    import piso_env_pkg::*;

    // Include config (not in a sub-package due to wide usage)
    `include "config/piso_config.sv"
endpackage