package piso_agent_pkg;
    import uvm_pkg::*;
    import piso_pkg::piso_config;
    import piso_sequences_pkg::piso_seq_item;
    `include "uvm_macros.svh"

    `include "piso_driver.sv"
    `include "piso_monitor.sv"
    `include "piso_sequencer.sv"
    `include "piso_agent.sv"
endpackage