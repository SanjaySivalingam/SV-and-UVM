package piso_env_pkg;
    import uvm_pkg::*;
    import piso_sequences_pkg::*;
    import piso_agent_pkg::*;
    `include "uvm_macros.svh"

    `include "piso_scoreboard.sv"
    `include "piso_coverage.sv"
    `include "piso_virtual_sequencer.sv"
    `include "piso_env.sv"
endpackage